`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Joshua Horwitz
// Create Date: 04/16/2015 10:04:05 PM
// 
//////////////////////////////////////////////////////////////////////////////////


module memory_mapper(
    input [1:0] unit_select,
    input [31:0] keyboard,
    input [31:0] screen,
    input [31:0] data_mem,
    output [31:0] to_mips
    );
    
    
    
endmodule
